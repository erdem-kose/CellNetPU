LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mpu IS
PORT (
	zio : INOUT STD_LOGIC;
	rzq : INOUT STD_LOGIC;
	mcbx_dram_we_n : OUT STD_LOGIC;
	mcbx_dram_udqs_n : INOUT STD_LOGIC;
	mcbx_dram_udqs : INOUT STD_LOGIC;
	mcbx_dram_udm : OUT STD_LOGIC;
	mcbx_dram_ras_n : OUT STD_LOGIC;
	mcbx_dram_odt : OUT STD_LOGIC;
	mcbx_dram_ldm : OUT STD_LOGIC;
	mcbx_dram_dqs_n : INOUT STD_LOGIC;
	mcbx_dram_dqs : INOUT STD_LOGIC;
	mcbx_dram_dq : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	mcbx_dram_clk_n : OUT STD_LOGIC;
	mcbx_dram_clk : OUT STD_LOGIC;
	mcbx_dram_cke : OUT STD_LOGIC;
	mcbx_dram_cas_n : OUT STD_LOGIC;
	mcbx_dram_ba : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
	mcbx_dram_addr : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	RESET : IN STD_LOGIC;
	QSPI_FLASH_SS : INOUT STD_LOGIC;
	QSPI_FLASH_SCLK : INOUT STD_LOGIC;
	QSPI_FLASH_IO1 : INOUT STD_LOGIC;
	QSPI_FLASH_IO0 : INOUT STD_LOGIC;
	GCLK : IN STD_LOGIC;
	Ethernet_Lite_TX_EN : OUT STD_LOGIC;
	Ethernet_Lite_TX_CLK : IN STD_LOGIC;
	Ethernet_Lite_TXD : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	Ethernet_Lite_RX_ER : IN STD_LOGIC;
	Ethernet_Lite_RX_DV : IN STD_LOGIC;
	Ethernet_Lite_RX_CLK : IN STD_LOGIC;
	Ethernet_Lite_RXD : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	Ethernet_Lite_PHY_RST_N : OUT STD_LOGIC;
	Ethernet_Lite_MDIO : INOUT STD_LOGIC;
	Ethernet_Lite_MDC : OUT STD_LOGIC;
	Ethernet_Lite_CRS : IN STD_LOGIC;
	Ethernet_Lite_COL : IN STD_LOGIC;
	iomodule_0_UART_Rx : IN STD_LOGIC;
	iomodule_0_UART_Tx : OUT STD_LOGIC;
	iomodule_0_GPO1 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	iomodule_0_GPI1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_i : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_u00 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_u01 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_u02 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_u10 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_u12 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_u11 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_u20 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_u21 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_u22 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_x00 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_x02 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_x01 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_x11 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_x10 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_x12 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_x20 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_x22 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	error_x21 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	u_data_in : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	u_data_out : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	u_address : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
	u_we : OUT STD_LOGIC;
	x_data_in : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	x_data_out : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	x_address : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
	x_we : OUT STD_LOGIC;
	ideal_address : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
	ideal_we : OUT STD_LOGIC;
	ideal_data_in : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	ideal_data_out : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_A00 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_A01 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_A02 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_A10 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_A11 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_A12 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_A20 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_A21 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_A22 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_B00 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_B01 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_B02 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_B10 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_B11 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_B12 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_B20 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_B21 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_B22 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_I : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_xbnd : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	template_ubnd : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END mpu;

ARCHITECTURE STRUCTURE OF mpu IS

BEGIN
END ARCHITECTURE STRUCTURE;
